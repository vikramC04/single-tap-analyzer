/*****************************************************************************
 *                                                                           *
 * Module:       Lab5                                                       *
 * Description:                                                              *
 *      This module is the top level module of SE2DA4 Lab 5                    *
 *                                                                           *
 *****************************************************************************/

module lab5 (
input				CLOCK_50,			// DONE
input		[0:0]	KEY, 					// DONE (for reset)
input 	[7:0] SW,               // DONE
output 	[7:0] LEDR,					// DONE

// Bidirectionals
inout		[15:0]		DRAM_DQ,		// DONE

// Outputs
// These outputs were exported so we can signal tap them. The entire system is actually contained within the sopc_system controller module.
output		[12:0]	DRAM_ADDR,	// DONE
output 		[1:0]		DRAM_BA,		// DONE
output					DRAM_LDQM,  // DONE data mask; when it is low, the DQ is valid for reading and writing. 
output					DRAM_UDQM,	// DONE
output					DRAM_RAS_N,	// DONE
output 					DRAM_CAS_N,	// DONE
output 					DRAM_CLK,	// DONE
output					DRAM_CKE,	// DONE
output 					DRAM_WE_N,	// DONE
output 					DRAM_CS_N	// DONE
);


// Internal Wires

assign LEDR=SW;

// Instantiate your sopc_system module generated by Platform Designer. (This refers to the system that we will be generating using the Platform designer.
// The SDRAM_Controller.v will be turned into a custom component which we will connect to the processor. This entire system is than instantiated below).

sopc_system  controller (
		.clk_clk(CLOCK_50),					// clk.clk
		.reset_reset_n(KEY[0]),				// reset.reset_n
		.sdram_addr_address(DRAM_ADDR),
		.sdram_ba_readdata(DRAM_BA),
		.sdram_cas_n_writeresponsevalid_n(DRAM_CAS_N),
		.sdram_cke_writeresponsevalid_n(DRAM_CKE),
		.sdram_clk_clk(DRAM_CLK),
		.sdram_cs_n_writeresponsevalid_n(DRAM_CS_N),
		.sdram_dq_export(DRAM_DQ),
		.sdram_ldqm_writeresponsevalid_n(DRAM_LDQM),
		.sdram_ras_n_writeresponsevalid_n(DRAM_RAS_N),
		.sdram_udqm_writeresponsevalid_n(DRAM_UDQM),
		.sdram_we_n_writeresponsevalid_n(DRAM_WE_N)
	);
	
endmodule
